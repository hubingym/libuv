module main

import libuv

fn main() {
    println('hello world')
}
